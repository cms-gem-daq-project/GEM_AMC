------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity trigger is
    generic(
        g_NUM_OF_OHs        : integer;
        g_NUM_TRIG_TX_LINKS : integer;
        g_USE_TRIG_TX_LINKS : boolean
    );
    port(
        -- reset
        reset_i             : in  std_logic;
        
        -- TTC
        ttc_clk_i           : in  t_ttc_clks;
        ttc_cmds_i          : in  t_ttc_cmds;

        -- Sbit cluster inputs
        sbit_clusters_i     : in t_oh_sbits_arr(g_NUM_OF_OHs - 1 downto 0);
        sbit_link_status_i  : in t_oh_sbit_links_arr(g_NUM_OF_OHs - 1 downto 0);

        -- Outputs
        trig_led_o          : out std_logic;
        trig_tx_data_arr_o  : out t_std234_array(g_NUM_TRIG_TX_LINKS - 1 downto 0);

        -- IPbus
        ipb_reset_i         : in  std_logic;
        ipb_clk_i           : in  std_logic;
        ipb_miso_o          : out ipb_rbus;
        ipb_mosi_i          : in  ipb_wbus
    );
end trigger;

architecture trigger_arch of trigger is
    
    signal reset_global         : std_logic;
    signal reset_local          : std_logic;
    signal reset                : std_logic;
    signal reset_cnt            : std_logic;
    
    signal oh_mask              : std_logic_vector(23 downto 0) := (others => '0');
    signal oh_triggers          : std_logic_vector(g_NUM_OF_OHs - 1 downto 0) := (others => '0');
    signal oh_num_valid_arr     : t_std4_array(g_NUM_OF_OHs - 1 downto 0);
    signal or_trigger           : std_logic;
        
    signal sbitmon_reset        : std_logic;
    signal sbitmon_sbits        : t_oh_sbits;
    signal sbitmon_l1a_delay    : std_logic_vector(31 downto 0);
    signal sbitmon_link_select  : std_logic_vector(3 downto 0);
    
    -- counters
    signal or_trigger_rate      : std_logic_vector(31 downto 0); 
    signal or_trigger_cnt       : std_logic_vector(31 downto 0); 
    
    -- OH counters
    signal sbit_overflow_cnt    : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal missed_comma_cnt     : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal link_overflow_cnt    : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal link_underflow_cnt   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal sync_word_cnt        : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trigger_rate         : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trigger_cnt          : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal cluster_cnt_rate     : t_std32_array((g_NUM_OF_OHs * 9) - 1 downto 0);
    signal cluster_cnt          : t_std32_array((g_NUM_OF_OHs * 9) - 1 downto 0);

    -- trigger output to EMTF
    signal sector_id            : std_logic_vector(3 downto 0);
    
    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------
    
begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clk_i.clk_40,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;

    --== Trigger ==--
    
    or_trigger <= or_reduce(oh_triggers);

    i_or_trigger_rate : entity work.rate_counter
        generic map(
            g_CLK_FREQUENCY => C_TTC_CLK_FREQUENCY_SLV,
            g_COUNTER_WIDTH => 32
        )
        port map(
            clk_i   => ttc_clk_i.clk_40,
            reset_i => reset or reset_cnt,
            en_i    => or_trigger,
            rate_o  => or_trigger_rate
        );

    i_or_trigger_cnt: entity work.counter
        generic map(
            g_COUNTER_WIDTH  => 32,
            g_ALLOW_ROLLOVER => FALSE
        )
        port map(
            ref_clk_i => ttc_clk_i.clk_40,
            reset_i   => reset or reset_cnt,
            en_i      => or_trigger,
            count_o   => or_trigger_cnt
        );
    
    i_led_pulse : entity work.pulse_extend
        generic map(
            DELAY_CNT_LENGTH => C_LED_PULSE_LENGTH_TTC_CLK'length
        )
        port map(
            clk_i          => ttc_clk_i.clk_40,
            rst_i          => reset,
            pulse_length_i => C_LED_PULSE_LENGTH_TTC_CLK,
            pulse_i        => or_trigger,
            pulse_o        => trig_led_o
        );
    
    --== Links ==--
        
    -- TODO: imlpement link synchronization by looking for sync words after each resync and delay the data of all links to match the latest one (use FIFOs for that) 
    g_input_processors:
    for i in 0 to g_NUM_OF_OHs - 1 generate
        
        i_input_processor: entity work.trigger_input_processor
            port map(
                reset_i              => reset,
                reset_cnt_i          => reset_cnt,
                clk_i                => ttc_clk_i.clk_40,
                sbit_clusters_i      => sbit_clusters_i(i),
                link_status_i        => sbit_link_status_i(i),
                masked_i             => oh_mask(i),
                trigger_o            => oh_triggers(i),
                num_valid_clusters_o => oh_num_valid_arr(i),
                sbit_overflow_cnt_o  => sbit_overflow_cnt(i),
                missed_comma_cnt_o   => missed_comma_cnt(i),
                link_overflow_cnt_o  => link_overflow_cnt(i),
                link_underflow_cnt_o => link_underflow_cnt(i),
                sync_word_cnt_o      => sync_word_cnt(i),
                cluster_cnt_rate_o   => cluster_cnt_rate(((i + 1) * 9) - 1 downto i * 9),
                trigger_rate_o       => trigger_rate(i),
                cluster_cnt_o        => cluster_cnt(((i + 1) * 9) - 1 downto i * 9),
                trigger_cnt_o        => trigger_cnt(i)
            );
        
    end generate;

    --== SBit monitor ==--
    
    i_sbit_monitor : entity work.sbit_monitor
        generic map(
            g_NUM_OF_OHs => g_NUM_OF_OHs
        )
        port map(
            reset_i         => sbitmon_reset,
            ttc_clk_i       => ttc_clk_i,
            ttc_cmds_i      => ttc_cmds_i,
            link_select_i   => sbitmon_link_select,
            sbit_clusters_i => sbit_clusters_i,
            sbit_trigger_i  => oh_triggers,
            frozen_sbits_o  => sbitmon_sbits,
            l1a_dealy_o     => sbitmon_l1a_delay
        );
    
    --== Output ==--
    
    g_use_trig_out : if g_USE_TRIG_TX_LINKS generate
        i_trig_output : entity work.trigger_output
            generic map(
                g_NUM_OF_OHs        => g_NUM_OF_OHs,
                g_NUM_TRIG_TX_LINKS => g_NUM_TRIG_TX_LINKS
            )
            port map(
                reset_i            => reset_i,
                ttc_clk_i          => ttc_clk_i,
                ttc_cmds_i         => ttc_cmds_i,
                sbit_clusters_i    => sbit_clusters_i,
                sbit_num_valid_i   => oh_num_valid_arr,
                oh_triggers_i      => oh_triggers,
                oh_mask_i          => oh_mask(g_NUM_OF_OHs - 1 downto 0),
                sbit_link_status_i => sbit_link_status_i,
                sector_id_i        => sector_id,
                trig_tx_data_arr_o => trig_tx_data_arr_o
            );
    end generate;

    g_fake_trig_out : if not g_USE_TRIG_TX_LINKS generate
        g_fake_trig_link : for i in 0 to g_NUM_TRIG_TX_LINKS - 1 generate
            trig_tx_data_arr_o(i) <= (others => '1');
        end generate;
    end generate;    
    
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_TRIGGER_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_TRIGGER_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_TRIGGER_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => ttc_clk_i.clk_40,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"000";
    regs_addresses(1)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"001";
    regs_addresses(2)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"002";
    regs_addresses(3)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"010";
    regs_addresses(4)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"011";
    regs_addresses(5)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"080";
    regs_addresses(6)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"081";
    regs_addresses(7)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"082";
    regs_addresses(8)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"083";
    regs_addresses(9)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"084";
    regs_addresses(10)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"085";
    regs_addresses(11)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"086";
    regs_addresses(12)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"087";
    regs_addresses(13)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"088";
    regs_addresses(14)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"089";
    regs_addresses(15)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"08a";
    regs_addresses(16)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"100";
    regs_addresses(17)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"101";
    regs_addresses(18)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"110";
    regs_addresses(19)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"111";
    regs_addresses(20)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"112";
    regs_addresses(21)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"113";
    regs_addresses(22)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"114";
    regs_addresses(23)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"115";
    regs_addresses(24)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"116";
    regs_addresses(25)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"117";
    regs_addresses(26)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"118";
    regs_addresses(27)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"120";
    regs_addresses(28)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"121";
    regs_addresses(29)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"122";
    regs_addresses(30)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"123";
    regs_addresses(31)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"124";
    regs_addresses(32)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"125";
    regs_addresses(33)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"126";
    regs_addresses(34)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"127";
    regs_addresses(35)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"128";
    regs_addresses(36)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a0";
    regs_addresses(37)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a1";
    regs_addresses(38)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a3";
    regs_addresses(39)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a4";
    regs_addresses(40)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a5";
    regs_addresses(41)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"200";
    regs_addresses(42)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"201";
    regs_addresses(43)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"210";
    regs_addresses(44)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"211";
    regs_addresses(45)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"212";
    regs_addresses(46)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"213";
    regs_addresses(47)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"214";
    regs_addresses(48)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"215";
    regs_addresses(49)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"216";
    regs_addresses(50)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"217";
    regs_addresses(51)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"218";
    regs_addresses(52)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"220";
    regs_addresses(53)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"221";
    regs_addresses(54)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"222";
    regs_addresses(55)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"223";
    regs_addresses(56)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"224";
    regs_addresses(57)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"225";
    regs_addresses(58)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"226";
    regs_addresses(59)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"227";
    regs_addresses(60)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"228";
    regs_addresses(61)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a0";
    regs_addresses(62)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a1";
    regs_addresses(63)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a3";
    regs_addresses(64)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a4";
    regs_addresses(65)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a5";
    regs_addresses(66)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"300";
    regs_addresses(67)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"301";
    regs_addresses(68)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"310";
    regs_addresses(69)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"311";
    regs_addresses(70)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"312";
    regs_addresses(71)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"313";
    regs_addresses(72)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"314";
    regs_addresses(73)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"315";
    regs_addresses(74)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"316";
    regs_addresses(75)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"317";
    regs_addresses(76)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"318";
    regs_addresses(77)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"320";
    regs_addresses(78)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"321";
    regs_addresses(79)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"322";
    regs_addresses(80)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"323";
    regs_addresses(81)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"324";
    regs_addresses(82)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"325";
    regs_addresses(83)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"326";
    regs_addresses(84)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"327";
    regs_addresses(85)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"328";
    regs_addresses(86)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"3a0";
    regs_addresses(87)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"3a1";
    regs_addresses(88)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"3a3";
    regs_addresses(89)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"3a4";
    regs_addresses(90)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"3a5";
    regs_addresses(91)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"400";
    regs_addresses(92)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"401";
    regs_addresses(93)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"410";
    regs_addresses(94)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"411";
    regs_addresses(95)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"412";
    regs_addresses(96)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"413";
    regs_addresses(97)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"414";
    regs_addresses(98)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"415";
    regs_addresses(99)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"416";
    regs_addresses(100)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"417";
    regs_addresses(101)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"418";
    regs_addresses(102)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"420";
    regs_addresses(103)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"421";
    regs_addresses(104)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"422";
    regs_addresses(105)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"423";
    regs_addresses(106)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"424";
    regs_addresses(107)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"425";
    regs_addresses(108)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"426";
    regs_addresses(109)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"427";
    regs_addresses(110)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"428";
    regs_addresses(111)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"4a0";
    regs_addresses(112)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"4a1";
    regs_addresses(113)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"4a3";
    regs_addresses(114)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"4a4";
    regs_addresses(115)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"4a5";
    regs_addresses(116)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"500";
    regs_addresses(117)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"501";
    regs_addresses(118)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"510";
    regs_addresses(119)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"511";
    regs_addresses(120)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"512";
    regs_addresses(121)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"513";
    regs_addresses(122)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"514";
    regs_addresses(123)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"515";
    regs_addresses(124)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"516";
    regs_addresses(125)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"517";
    regs_addresses(126)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"518";
    regs_addresses(127)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"520";
    regs_addresses(128)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"521";
    regs_addresses(129)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"522";
    regs_addresses(130)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"523";
    regs_addresses(131)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"524";
    regs_addresses(132)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"525";
    regs_addresses(133)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"526";
    regs_addresses(134)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"527";
    regs_addresses(135)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"528";
    regs_addresses(136)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"5a0";
    regs_addresses(137)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"5a1";
    regs_addresses(138)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"5a3";
    regs_addresses(139)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"5a4";
    regs_addresses(140)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"5a5";
    regs_addresses(141)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"600";
    regs_addresses(142)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"601";
    regs_addresses(143)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"610";
    regs_addresses(144)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"611";
    regs_addresses(145)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"612";
    regs_addresses(146)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"613";
    regs_addresses(147)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"614";
    regs_addresses(148)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"615";
    regs_addresses(149)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"616";
    regs_addresses(150)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"617";
    regs_addresses(151)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"618";
    regs_addresses(152)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"620";
    regs_addresses(153)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"621";
    regs_addresses(154)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"622";
    regs_addresses(155)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"623";
    regs_addresses(156)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"624";
    regs_addresses(157)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"625";
    regs_addresses(158)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"626";
    regs_addresses(159)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"627";
    regs_addresses(160)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"628";
    regs_addresses(161)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"6a0";
    regs_addresses(162)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"6a1";
    regs_addresses(163)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"6a3";
    regs_addresses(164)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"6a4";
    regs_addresses(165)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"6a5";
    regs_addresses(166)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"700";
    regs_addresses(167)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"701";
    regs_addresses(168)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"710";
    regs_addresses(169)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"711";
    regs_addresses(170)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"712";
    regs_addresses(171)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"713";
    regs_addresses(172)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"714";
    regs_addresses(173)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"715";
    regs_addresses(174)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"716";
    regs_addresses(175)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"717";
    regs_addresses(176)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"718";
    regs_addresses(177)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"720";
    regs_addresses(178)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"721";
    regs_addresses(179)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"722";
    regs_addresses(180)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"723";
    regs_addresses(181)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"724";
    regs_addresses(182)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"725";
    regs_addresses(183)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"726";
    regs_addresses(184)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"727";
    regs_addresses(185)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"728";
    regs_addresses(186)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"7a0";
    regs_addresses(187)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"7a1";
    regs_addresses(188)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"7a3";
    regs_addresses(189)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"7a4";
    regs_addresses(190)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"7a5";
    regs_addresses(191)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"800";
    regs_addresses(192)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"801";
    regs_addresses(193)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"810";
    regs_addresses(194)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"811";
    regs_addresses(195)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"812";
    regs_addresses(196)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"813";
    regs_addresses(197)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"814";
    regs_addresses(198)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"815";
    regs_addresses(199)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"816";
    regs_addresses(200)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"817";
    regs_addresses(201)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"818";
    regs_addresses(202)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"820";
    regs_addresses(203)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"821";
    regs_addresses(204)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"822";
    regs_addresses(205)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"823";
    regs_addresses(206)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"824";
    regs_addresses(207)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"825";
    regs_addresses(208)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"826";
    regs_addresses(209)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"827";
    regs_addresses(210)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"828";
    regs_addresses(211)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"8a0";
    regs_addresses(212)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"8a1";
    regs_addresses(213)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"8a3";
    regs_addresses(214)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"8a4";
    regs_addresses(215)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"8a5";
    regs_addresses(216)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"900";
    regs_addresses(217)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"901";
    regs_addresses(218)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"910";
    regs_addresses(219)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"911";
    regs_addresses(220)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"912";
    regs_addresses(221)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"913";
    regs_addresses(222)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"914";
    regs_addresses(223)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"915";
    regs_addresses(224)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"916";
    regs_addresses(225)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"917";
    regs_addresses(226)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"918";
    regs_addresses(227)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"920";
    regs_addresses(228)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"921";
    regs_addresses(229)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"922";
    regs_addresses(230)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"923";
    regs_addresses(231)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"924";
    regs_addresses(232)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"925";
    regs_addresses(233)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"926";
    regs_addresses(234)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"927";
    regs_addresses(235)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"928";
    regs_addresses(236)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"9a0";
    regs_addresses(237)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"9a1";
    regs_addresses(238)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"9a3";
    regs_addresses(239)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"9a4";
    regs_addresses(240)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"9a5";
    regs_addresses(241)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a00";
    regs_addresses(242)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a01";
    regs_addresses(243)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a10";
    regs_addresses(244)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a11";
    regs_addresses(245)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a12";
    regs_addresses(246)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a13";
    regs_addresses(247)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a14";
    regs_addresses(248)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a15";
    regs_addresses(249)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a16";
    regs_addresses(250)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a17";
    regs_addresses(251)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a18";
    regs_addresses(252)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a20";
    regs_addresses(253)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a21";
    regs_addresses(254)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a22";
    regs_addresses(255)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a23";
    regs_addresses(256)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a24";
    regs_addresses(257)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a25";
    regs_addresses(258)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a26";
    regs_addresses(259)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a27";
    regs_addresses(260)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"a28";
    regs_addresses(261)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"aa0";
    regs_addresses(262)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"aa1";
    regs_addresses(263)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"aa3";
    regs_addresses(264)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"aa4";
    regs_addresses(265)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"aa5";
    regs_addresses(266)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b00";
    regs_addresses(267)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b01";
    regs_addresses(268)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b10";
    regs_addresses(269)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b11";
    regs_addresses(270)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b12";
    regs_addresses(271)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b13";
    regs_addresses(272)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b14";
    regs_addresses(273)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b15";
    regs_addresses(274)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b16";
    regs_addresses(275)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b17";
    regs_addresses(276)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b18";
    regs_addresses(277)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b20";
    regs_addresses(278)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b21";
    regs_addresses(279)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b22";
    regs_addresses(280)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b23";
    regs_addresses(281)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b24";
    regs_addresses(282)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b25";
    regs_addresses(283)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b26";
    regs_addresses(284)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b27";
    regs_addresses(285)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"b28";
    regs_addresses(286)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ba0";
    regs_addresses(287)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ba1";
    regs_addresses(288)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ba3";
    regs_addresses(289)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ba4";
    regs_addresses(290)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ba5";
    regs_addresses(291)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c00";
    regs_addresses(292)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c01";
    regs_addresses(293)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c10";
    regs_addresses(294)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c11";
    regs_addresses(295)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c12";
    regs_addresses(296)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c13";
    regs_addresses(297)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c14";
    regs_addresses(298)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c15";
    regs_addresses(299)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c16";
    regs_addresses(300)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c17";
    regs_addresses(301)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c18";
    regs_addresses(302)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c20";
    regs_addresses(303)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c21";
    regs_addresses(304)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c22";
    regs_addresses(305)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c23";
    regs_addresses(306)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c24";
    regs_addresses(307)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c25";
    regs_addresses(308)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c26";
    regs_addresses(309)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c27";
    regs_addresses(310)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"c28";
    regs_addresses(311)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ca0";
    regs_addresses(312)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ca1";
    regs_addresses(313)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ca3";
    regs_addresses(314)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ca4";
    regs_addresses(315)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"ca5";

    -- Connect read signals
    regs_read_arr(2)(REG_TRIGGER_CTRL_OH_KILL_MASK_MSB downto REG_TRIGGER_CTRL_OH_KILL_MASK_LSB) <= oh_mask;
    regs_read_arr(2)(REG_TRIGGER_CTRL_SECTOR_ID_MSB downto REG_TRIGGER_CTRL_SECTOR_ID_LSB) <= sector_id;
    regs_read_arr(3)(REG_TRIGGER_STATUS_OR_TRIGGER_RATE_MSB downto REG_TRIGGER_STATUS_OR_TRIGGER_RATE_LSB) <= or_trigger_rate;
    regs_read_arr(4)(REG_TRIGGER_STATUS_OR_TRIGGER_CNT_MSB downto REG_TRIGGER_STATUS_OR_TRIGGER_CNT_LSB) <= or_trigger_cnt;
    regs_read_arr(6)(REG_TRIGGER_SBIT_MONITOR_OH_SELECT_MSB downto REG_TRIGGER_SBIT_MONITOR_OH_SELECT_LSB) <= sbitmon_link_select;
    regs_read_arr(7)(REG_TRIGGER_SBIT_MONITOR_CLUSTER0_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER0_LSB) <= '0' & sbitmon_sbits(0).size & '0' & sbitmon_sbits(0).address;
    regs_read_arr(8)(REG_TRIGGER_SBIT_MONITOR_CLUSTER1_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER1_LSB) <= '0' & sbitmon_sbits(1).size & '0' & sbitmon_sbits(1).address;
    regs_read_arr(9)(REG_TRIGGER_SBIT_MONITOR_CLUSTER2_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER2_LSB) <= '0' & sbitmon_sbits(2).size & '0' & sbitmon_sbits(2).address;
    regs_read_arr(10)(REG_TRIGGER_SBIT_MONITOR_CLUSTER3_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER3_LSB) <= '0' & sbitmon_sbits(3).size & '0' & sbitmon_sbits(3).address;
    regs_read_arr(11)(REG_TRIGGER_SBIT_MONITOR_CLUSTER4_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER4_LSB) <= '0' & sbitmon_sbits(4).size & '0' & sbitmon_sbits(4).address;
    regs_read_arr(12)(REG_TRIGGER_SBIT_MONITOR_CLUSTER5_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER5_LSB) <= '0' & sbitmon_sbits(5).size & '0' & sbitmon_sbits(5).address;
    regs_read_arr(13)(REG_TRIGGER_SBIT_MONITOR_CLUSTER6_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER6_LSB) <= '0' & sbitmon_sbits(6).size & '0' & sbitmon_sbits(6).address;
    regs_read_arr(14)(REG_TRIGGER_SBIT_MONITOR_CLUSTER7_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER7_LSB) <= '0' & sbitmon_sbits(7).size & '0' & sbitmon_sbits(7).address;
    regs_read_arr(15)(REG_TRIGGER_SBIT_MONITOR_L1A_DELAY_MSB downto REG_TRIGGER_SBIT_MONITOR_L1A_DELAY_LSB) <= sbitmon_l1a_delay;
    regs_read_arr(16)(REG_TRIGGER_OH0_TRIGGER_RATE_MSB downto REG_TRIGGER_OH0_TRIGGER_RATE_LSB) <= trigger_rate(0);
    regs_read_arr(17)(REG_TRIGGER_OH0_TRIGGER_CNT_MSB downto REG_TRIGGER_OH0_TRIGGER_CNT_LSB) <= trigger_cnt(0);
    regs_read_arr(18)(REG_TRIGGER_OH0_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 0);
    regs_read_arr(19)(REG_TRIGGER_OH0_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 1);
    regs_read_arr(20)(REG_TRIGGER_OH0_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 2);
    regs_read_arr(21)(REG_TRIGGER_OH0_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 3);
    regs_read_arr(22)(REG_TRIGGER_OH0_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 4);
    regs_read_arr(23)(REG_TRIGGER_OH0_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 5);
    regs_read_arr(24)(REG_TRIGGER_OH0_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 6);
    regs_read_arr(25)(REG_TRIGGER_OH0_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 7);
    regs_read_arr(26)(REG_TRIGGER_OH0_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 8);
    regs_read_arr(27)(REG_TRIGGER_OH0_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(0 * 9 + 0);
    regs_read_arr(28)(REG_TRIGGER_OH0_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(0 * 9 + 1);
    regs_read_arr(29)(REG_TRIGGER_OH0_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(0 * 9 + 2);
    regs_read_arr(30)(REG_TRIGGER_OH0_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(0 * 9 + 3);
    regs_read_arr(31)(REG_TRIGGER_OH0_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(0 * 9 + 4);
    regs_read_arr(32)(REG_TRIGGER_OH0_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(0 * 9 + 5);
    regs_read_arr(33)(REG_TRIGGER_OH0_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(0 * 9 + 6);
    regs_read_arr(34)(REG_TRIGGER_OH0_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(0 * 9 + 7);
    regs_read_arr(35)(REG_TRIGGER_OH0_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(0 * 9 + 8);
    regs_read_arr(36)(REG_TRIGGER_OH0_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(0)(15 downto 0);
    regs_read_arr(36)(REG_TRIGGER_OH0_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(0)(31 downto 16);
    regs_read_arr(37)(REG_TRIGGER_OH0_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH0_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(0)(15 downto 0);
    regs_read_arr(37)(REG_TRIGGER_OH0_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH0_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(0)(31 downto 16);
    regs_read_arr(38)(REG_TRIGGER_OH0_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(0)(15 downto 0);
    regs_read_arr(38)(REG_TRIGGER_OH0_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(0)(31 downto 16);
    regs_read_arr(39)(REG_TRIGGER_OH0_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(0)(15 downto 0);
    regs_read_arr(39)(REG_TRIGGER_OH0_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(0)(31 downto 16);
    regs_read_arr(40)(REG_TRIGGER_OH0_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH0_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(0)(15 downto 0);
    regs_read_arr(40)(REG_TRIGGER_OH0_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH0_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(0)(31 downto 16);
    regs_read_arr(41)(REG_TRIGGER_OH1_TRIGGER_RATE_MSB downto REG_TRIGGER_OH1_TRIGGER_RATE_LSB) <= trigger_rate(1);
    regs_read_arr(42)(REG_TRIGGER_OH1_TRIGGER_CNT_MSB downto REG_TRIGGER_OH1_TRIGGER_CNT_LSB) <= trigger_cnt(1);
    regs_read_arr(43)(REG_TRIGGER_OH1_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 0);
    regs_read_arr(44)(REG_TRIGGER_OH1_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 1);
    regs_read_arr(45)(REG_TRIGGER_OH1_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 2);
    regs_read_arr(46)(REG_TRIGGER_OH1_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 3);
    regs_read_arr(47)(REG_TRIGGER_OH1_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 4);
    regs_read_arr(48)(REG_TRIGGER_OH1_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 5);
    regs_read_arr(49)(REG_TRIGGER_OH1_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 6);
    regs_read_arr(50)(REG_TRIGGER_OH1_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 7);
    regs_read_arr(51)(REG_TRIGGER_OH1_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 8);
    regs_read_arr(52)(REG_TRIGGER_OH1_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(1 * 9 + 0);
    regs_read_arr(53)(REG_TRIGGER_OH1_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(1 * 9 + 1);
    regs_read_arr(54)(REG_TRIGGER_OH1_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(1 * 9 + 2);
    regs_read_arr(55)(REG_TRIGGER_OH1_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(1 * 9 + 3);
    regs_read_arr(56)(REG_TRIGGER_OH1_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(1 * 9 + 4);
    regs_read_arr(57)(REG_TRIGGER_OH1_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(1 * 9 + 5);
    regs_read_arr(58)(REG_TRIGGER_OH1_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(1 * 9 + 6);
    regs_read_arr(59)(REG_TRIGGER_OH1_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(1 * 9 + 7);
    regs_read_arr(60)(REG_TRIGGER_OH1_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(1 * 9 + 8);
    regs_read_arr(61)(REG_TRIGGER_OH1_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(1)(15 downto 0);
    regs_read_arr(61)(REG_TRIGGER_OH1_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(1)(31 downto 16);
    regs_read_arr(62)(REG_TRIGGER_OH1_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH1_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(1)(15 downto 0);
    regs_read_arr(62)(REG_TRIGGER_OH1_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH1_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(1)(31 downto 16);
    regs_read_arr(63)(REG_TRIGGER_OH1_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(1)(15 downto 0);
    regs_read_arr(63)(REG_TRIGGER_OH1_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(1)(31 downto 16);
    regs_read_arr(64)(REG_TRIGGER_OH1_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(1)(15 downto 0);
    regs_read_arr(64)(REG_TRIGGER_OH1_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(1)(31 downto 16);
    regs_read_arr(65)(REG_TRIGGER_OH1_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH1_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(1)(15 downto 0);
    regs_read_arr(65)(REG_TRIGGER_OH1_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH1_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(1)(31 downto 16);
    regs_read_arr(66)(REG_TRIGGER_OH2_TRIGGER_RATE_MSB downto REG_TRIGGER_OH2_TRIGGER_RATE_LSB) <= trigger_rate(2);
    regs_read_arr(67)(REG_TRIGGER_OH2_TRIGGER_CNT_MSB downto REG_TRIGGER_OH2_TRIGGER_CNT_LSB) <= trigger_cnt(2);
    regs_read_arr(68)(REG_TRIGGER_OH2_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 0);
    regs_read_arr(69)(REG_TRIGGER_OH2_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 1);
    regs_read_arr(70)(REG_TRIGGER_OH2_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 2);
    regs_read_arr(71)(REG_TRIGGER_OH2_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 3);
    regs_read_arr(72)(REG_TRIGGER_OH2_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 4);
    regs_read_arr(73)(REG_TRIGGER_OH2_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 5);
    regs_read_arr(74)(REG_TRIGGER_OH2_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 6);
    regs_read_arr(75)(REG_TRIGGER_OH2_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 7);
    regs_read_arr(76)(REG_TRIGGER_OH2_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(2 * 9 + 8);
    regs_read_arr(77)(REG_TRIGGER_OH2_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(2 * 9 + 0);
    regs_read_arr(78)(REG_TRIGGER_OH2_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(2 * 9 + 1);
    regs_read_arr(79)(REG_TRIGGER_OH2_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(2 * 9 + 2);
    regs_read_arr(80)(REG_TRIGGER_OH2_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(2 * 9 + 3);
    regs_read_arr(81)(REG_TRIGGER_OH2_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(2 * 9 + 4);
    regs_read_arr(82)(REG_TRIGGER_OH2_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(2 * 9 + 5);
    regs_read_arr(83)(REG_TRIGGER_OH2_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(2 * 9 + 6);
    regs_read_arr(84)(REG_TRIGGER_OH2_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(2 * 9 + 7);
    regs_read_arr(85)(REG_TRIGGER_OH2_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH2_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(2 * 9 + 8);
    regs_read_arr(86)(REG_TRIGGER_OH2_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH2_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(2)(15 downto 0);
    regs_read_arr(86)(REG_TRIGGER_OH2_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH2_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(2)(31 downto 16);
    regs_read_arr(87)(REG_TRIGGER_OH2_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH2_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(2)(15 downto 0);
    regs_read_arr(87)(REG_TRIGGER_OH2_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH2_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(2)(31 downto 16);
    regs_read_arr(88)(REG_TRIGGER_OH2_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH2_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(2)(15 downto 0);
    regs_read_arr(88)(REG_TRIGGER_OH2_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH2_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(2)(31 downto 16);
    regs_read_arr(89)(REG_TRIGGER_OH2_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH2_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(2)(15 downto 0);
    regs_read_arr(89)(REG_TRIGGER_OH2_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH2_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(2)(31 downto 16);
    regs_read_arr(90)(REG_TRIGGER_OH2_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH2_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(2)(15 downto 0);
    regs_read_arr(90)(REG_TRIGGER_OH2_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH2_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(2)(31 downto 16);
    regs_read_arr(91)(REG_TRIGGER_OH3_TRIGGER_RATE_MSB downto REG_TRIGGER_OH3_TRIGGER_RATE_LSB) <= trigger_rate(3);
    regs_read_arr(92)(REG_TRIGGER_OH3_TRIGGER_CNT_MSB downto REG_TRIGGER_OH3_TRIGGER_CNT_LSB) <= trigger_cnt(3);
    regs_read_arr(93)(REG_TRIGGER_OH3_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 0);
    regs_read_arr(94)(REG_TRIGGER_OH3_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 1);
    regs_read_arr(95)(REG_TRIGGER_OH3_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 2);
    regs_read_arr(96)(REG_TRIGGER_OH3_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 3);
    regs_read_arr(97)(REG_TRIGGER_OH3_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 4);
    regs_read_arr(98)(REG_TRIGGER_OH3_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 5);
    regs_read_arr(99)(REG_TRIGGER_OH3_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 6);
    regs_read_arr(100)(REG_TRIGGER_OH3_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 7);
    regs_read_arr(101)(REG_TRIGGER_OH3_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(3 * 9 + 8);
    regs_read_arr(102)(REG_TRIGGER_OH3_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(3 * 9 + 0);
    regs_read_arr(103)(REG_TRIGGER_OH3_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(3 * 9 + 1);
    regs_read_arr(104)(REG_TRIGGER_OH3_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(3 * 9 + 2);
    regs_read_arr(105)(REG_TRIGGER_OH3_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(3 * 9 + 3);
    regs_read_arr(106)(REG_TRIGGER_OH3_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(3 * 9 + 4);
    regs_read_arr(107)(REG_TRIGGER_OH3_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(3 * 9 + 5);
    regs_read_arr(108)(REG_TRIGGER_OH3_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(3 * 9 + 6);
    regs_read_arr(109)(REG_TRIGGER_OH3_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(3 * 9 + 7);
    regs_read_arr(110)(REG_TRIGGER_OH3_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH3_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(3 * 9 + 8);
    regs_read_arr(111)(REG_TRIGGER_OH3_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH3_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(3)(15 downto 0);
    regs_read_arr(111)(REG_TRIGGER_OH3_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH3_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(3)(31 downto 16);
    regs_read_arr(112)(REG_TRIGGER_OH3_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH3_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(3)(15 downto 0);
    regs_read_arr(112)(REG_TRIGGER_OH3_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH3_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(3)(31 downto 16);
    regs_read_arr(113)(REG_TRIGGER_OH3_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH3_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(3)(15 downto 0);
    regs_read_arr(113)(REG_TRIGGER_OH3_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH3_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(3)(31 downto 16);
    regs_read_arr(114)(REG_TRIGGER_OH3_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH3_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(3)(15 downto 0);
    regs_read_arr(114)(REG_TRIGGER_OH3_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH3_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(3)(31 downto 16);
    regs_read_arr(115)(REG_TRIGGER_OH3_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH3_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(3)(15 downto 0);
    regs_read_arr(115)(REG_TRIGGER_OH3_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH3_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(3)(31 downto 16);
    regs_read_arr(116)(REG_TRIGGER_OH4_TRIGGER_RATE_MSB downto REG_TRIGGER_OH4_TRIGGER_RATE_LSB) <= trigger_rate(4);
    regs_read_arr(117)(REG_TRIGGER_OH4_TRIGGER_CNT_MSB downto REG_TRIGGER_OH4_TRIGGER_CNT_LSB) <= trigger_cnt(4);
    regs_read_arr(118)(REG_TRIGGER_OH4_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 0);
    regs_read_arr(119)(REG_TRIGGER_OH4_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 1);
    regs_read_arr(120)(REG_TRIGGER_OH4_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 2);
    regs_read_arr(121)(REG_TRIGGER_OH4_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 3);
    regs_read_arr(122)(REG_TRIGGER_OH4_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 4);
    regs_read_arr(123)(REG_TRIGGER_OH4_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 5);
    regs_read_arr(124)(REG_TRIGGER_OH4_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 6);
    regs_read_arr(125)(REG_TRIGGER_OH4_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 7);
    regs_read_arr(126)(REG_TRIGGER_OH4_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(4 * 9 + 8);
    regs_read_arr(127)(REG_TRIGGER_OH4_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(4 * 9 + 0);
    regs_read_arr(128)(REG_TRIGGER_OH4_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(4 * 9 + 1);
    regs_read_arr(129)(REG_TRIGGER_OH4_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(4 * 9 + 2);
    regs_read_arr(130)(REG_TRIGGER_OH4_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(4 * 9 + 3);
    regs_read_arr(131)(REG_TRIGGER_OH4_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(4 * 9 + 4);
    regs_read_arr(132)(REG_TRIGGER_OH4_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(4 * 9 + 5);
    regs_read_arr(133)(REG_TRIGGER_OH4_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(4 * 9 + 6);
    regs_read_arr(134)(REG_TRIGGER_OH4_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(4 * 9 + 7);
    regs_read_arr(135)(REG_TRIGGER_OH4_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH4_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(4 * 9 + 8);
    regs_read_arr(136)(REG_TRIGGER_OH4_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH4_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(4)(15 downto 0);
    regs_read_arr(136)(REG_TRIGGER_OH4_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH4_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(4)(31 downto 16);
    regs_read_arr(137)(REG_TRIGGER_OH4_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH4_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(4)(15 downto 0);
    regs_read_arr(137)(REG_TRIGGER_OH4_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH4_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(4)(31 downto 16);
    regs_read_arr(138)(REG_TRIGGER_OH4_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH4_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(4)(15 downto 0);
    regs_read_arr(138)(REG_TRIGGER_OH4_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH4_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(4)(31 downto 16);
    regs_read_arr(139)(REG_TRIGGER_OH4_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH4_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(4)(15 downto 0);
    regs_read_arr(139)(REG_TRIGGER_OH4_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH4_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(4)(31 downto 16);
    regs_read_arr(140)(REG_TRIGGER_OH4_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH4_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(4)(15 downto 0);
    regs_read_arr(140)(REG_TRIGGER_OH4_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH4_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(4)(31 downto 16);
    regs_read_arr(141)(REG_TRIGGER_OH5_TRIGGER_RATE_MSB downto REG_TRIGGER_OH5_TRIGGER_RATE_LSB) <= trigger_rate(5);
    regs_read_arr(142)(REG_TRIGGER_OH5_TRIGGER_CNT_MSB downto REG_TRIGGER_OH5_TRIGGER_CNT_LSB) <= trigger_cnt(5);
    regs_read_arr(143)(REG_TRIGGER_OH5_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 0);
    regs_read_arr(144)(REG_TRIGGER_OH5_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 1);
    regs_read_arr(145)(REG_TRIGGER_OH5_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 2);
    regs_read_arr(146)(REG_TRIGGER_OH5_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 3);
    regs_read_arr(147)(REG_TRIGGER_OH5_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 4);
    regs_read_arr(148)(REG_TRIGGER_OH5_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 5);
    regs_read_arr(149)(REG_TRIGGER_OH5_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 6);
    regs_read_arr(150)(REG_TRIGGER_OH5_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 7);
    regs_read_arr(151)(REG_TRIGGER_OH5_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(5 * 9 + 8);
    regs_read_arr(152)(REG_TRIGGER_OH5_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(5 * 9 + 0);
    regs_read_arr(153)(REG_TRIGGER_OH5_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(5 * 9 + 1);
    regs_read_arr(154)(REG_TRIGGER_OH5_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(5 * 9 + 2);
    regs_read_arr(155)(REG_TRIGGER_OH5_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(5 * 9 + 3);
    regs_read_arr(156)(REG_TRIGGER_OH5_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(5 * 9 + 4);
    regs_read_arr(157)(REG_TRIGGER_OH5_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(5 * 9 + 5);
    regs_read_arr(158)(REG_TRIGGER_OH5_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(5 * 9 + 6);
    regs_read_arr(159)(REG_TRIGGER_OH5_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(5 * 9 + 7);
    regs_read_arr(160)(REG_TRIGGER_OH5_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH5_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(5 * 9 + 8);
    regs_read_arr(161)(REG_TRIGGER_OH5_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH5_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(5)(15 downto 0);
    regs_read_arr(161)(REG_TRIGGER_OH5_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH5_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(5)(31 downto 16);
    regs_read_arr(162)(REG_TRIGGER_OH5_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH5_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(5)(15 downto 0);
    regs_read_arr(162)(REG_TRIGGER_OH5_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH5_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(5)(31 downto 16);
    regs_read_arr(163)(REG_TRIGGER_OH5_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH5_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(5)(15 downto 0);
    regs_read_arr(163)(REG_TRIGGER_OH5_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH5_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(5)(31 downto 16);
    regs_read_arr(164)(REG_TRIGGER_OH5_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH5_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(5)(15 downto 0);
    regs_read_arr(164)(REG_TRIGGER_OH5_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH5_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(5)(31 downto 16);
    regs_read_arr(165)(REG_TRIGGER_OH5_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH5_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(5)(15 downto 0);
    regs_read_arr(165)(REG_TRIGGER_OH5_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH5_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(5)(31 downto 16);
    regs_read_arr(166)(REG_TRIGGER_OH6_TRIGGER_RATE_MSB downto REG_TRIGGER_OH6_TRIGGER_RATE_LSB) <= trigger_rate(6);
    regs_read_arr(167)(REG_TRIGGER_OH6_TRIGGER_CNT_MSB downto REG_TRIGGER_OH6_TRIGGER_CNT_LSB) <= trigger_cnt(6);
    regs_read_arr(168)(REG_TRIGGER_OH6_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 0);
    regs_read_arr(169)(REG_TRIGGER_OH6_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 1);
    regs_read_arr(170)(REG_TRIGGER_OH6_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 2);
    regs_read_arr(171)(REG_TRIGGER_OH6_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 3);
    regs_read_arr(172)(REG_TRIGGER_OH6_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 4);
    regs_read_arr(173)(REG_TRIGGER_OH6_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 5);
    regs_read_arr(174)(REG_TRIGGER_OH6_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 6);
    regs_read_arr(175)(REG_TRIGGER_OH6_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 7);
    regs_read_arr(176)(REG_TRIGGER_OH6_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(6 * 9 + 8);
    regs_read_arr(177)(REG_TRIGGER_OH6_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(6 * 9 + 0);
    regs_read_arr(178)(REG_TRIGGER_OH6_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(6 * 9 + 1);
    regs_read_arr(179)(REG_TRIGGER_OH6_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(6 * 9 + 2);
    regs_read_arr(180)(REG_TRIGGER_OH6_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(6 * 9 + 3);
    regs_read_arr(181)(REG_TRIGGER_OH6_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(6 * 9 + 4);
    regs_read_arr(182)(REG_TRIGGER_OH6_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(6 * 9 + 5);
    regs_read_arr(183)(REG_TRIGGER_OH6_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(6 * 9 + 6);
    regs_read_arr(184)(REG_TRIGGER_OH6_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(6 * 9 + 7);
    regs_read_arr(185)(REG_TRIGGER_OH6_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH6_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(6 * 9 + 8);
    regs_read_arr(186)(REG_TRIGGER_OH6_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH6_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(6)(15 downto 0);
    regs_read_arr(186)(REG_TRIGGER_OH6_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH6_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(6)(31 downto 16);
    regs_read_arr(187)(REG_TRIGGER_OH6_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH6_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(6)(15 downto 0);
    regs_read_arr(187)(REG_TRIGGER_OH6_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH6_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(6)(31 downto 16);
    regs_read_arr(188)(REG_TRIGGER_OH6_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH6_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(6)(15 downto 0);
    regs_read_arr(188)(REG_TRIGGER_OH6_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH6_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(6)(31 downto 16);
    regs_read_arr(189)(REG_TRIGGER_OH6_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH6_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(6)(15 downto 0);
    regs_read_arr(189)(REG_TRIGGER_OH6_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH6_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(6)(31 downto 16);
    regs_read_arr(190)(REG_TRIGGER_OH6_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH6_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(6)(15 downto 0);
    regs_read_arr(190)(REG_TRIGGER_OH6_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH6_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(6)(31 downto 16);
    regs_read_arr(191)(REG_TRIGGER_OH7_TRIGGER_RATE_MSB downto REG_TRIGGER_OH7_TRIGGER_RATE_LSB) <= trigger_rate(7);
    regs_read_arr(192)(REG_TRIGGER_OH7_TRIGGER_CNT_MSB downto REG_TRIGGER_OH7_TRIGGER_CNT_LSB) <= trigger_cnt(7);
    regs_read_arr(193)(REG_TRIGGER_OH7_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 0);
    regs_read_arr(194)(REG_TRIGGER_OH7_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 1);
    regs_read_arr(195)(REG_TRIGGER_OH7_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 2);
    regs_read_arr(196)(REG_TRIGGER_OH7_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 3);
    regs_read_arr(197)(REG_TRIGGER_OH7_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 4);
    regs_read_arr(198)(REG_TRIGGER_OH7_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 5);
    regs_read_arr(199)(REG_TRIGGER_OH7_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 6);
    regs_read_arr(200)(REG_TRIGGER_OH7_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 7);
    regs_read_arr(201)(REG_TRIGGER_OH7_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(7 * 9 + 8);
    regs_read_arr(202)(REG_TRIGGER_OH7_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(7 * 9 + 0);
    regs_read_arr(203)(REG_TRIGGER_OH7_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(7 * 9 + 1);
    regs_read_arr(204)(REG_TRIGGER_OH7_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(7 * 9 + 2);
    regs_read_arr(205)(REG_TRIGGER_OH7_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(7 * 9 + 3);
    regs_read_arr(206)(REG_TRIGGER_OH7_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(7 * 9 + 4);
    regs_read_arr(207)(REG_TRIGGER_OH7_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(7 * 9 + 5);
    regs_read_arr(208)(REG_TRIGGER_OH7_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(7 * 9 + 6);
    regs_read_arr(209)(REG_TRIGGER_OH7_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(7 * 9 + 7);
    regs_read_arr(210)(REG_TRIGGER_OH7_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH7_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(7 * 9 + 8);
    regs_read_arr(211)(REG_TRIGGER_OH7_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH7_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(7)(15 downto 0);
    regs_read_arr(211)(REG_TRIGGER_OH7_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH7_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(7)(31 downto 16);
    regs_read_arr(212)(REG_TRIGGER_OH7_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH7_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(7)(15 downto 0);
    regs_read_arr(212)(REG_TRIGGER_OH7_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH7_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(7)(31 downto 16);
    regs_read_arr(213)(REG_TRIGGER_OH7_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH7_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(7)(15 downto 0);
    regs_read_arr(213)(REG_TRIGGER_OH7_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH7_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(7)(31 downto 16);
    regs_read_arr(214)(REG_TRIGGER_OH7_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH7_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(7)(15 downto 0);
    regs_read_arr(214)(REG_TRIGGER_OH7_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH7_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(7)(31 downto 16);
    regs_read_arr(215)(REG_TRIGGER_OH7_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH7_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(7)(15 downto 0);
    regs_read_arr(215)(REG_TRIGGER_OH7_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH7_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(7)(31 downto 16);
    regs_read_arr(216)(REG_TRIGGER_OH8_TRIGGER_RATE_MSB downto REG_TRIGGER_OH8_TRIGGER_RATE_LSB) <= trigger_rate(8);
    regs_read_arr(217)(REG_TRIGGER_OH8_TRIGGER_CNT_MSB downto REG_TRIGGER_OH8_TRIGGER_CNT_LSB) <= trigger_cnt(8);
    regs_read_arr(218)(REG_TRIGGER_OH8_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 0);
    regs_read_arr(219)(REG_TRIGGER_OH8_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 1);
    regs_read_arr(220)(REG_TRIGGER_OH8_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 2);
    regs_read_arr(221)(REG_TRIGGER_OH8_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 3);
    regs_read_arr(222)(REG_TRIGGER_OH8_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 4);
    regs_read_arr(223)(REG_TRIGGER_OH8_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 5);
    regs_read_arr(224)(REG_TRIGGER_OH8_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 6);
    regs_read_arr(225)(REG_TRIGGER_OH8_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 7);
    regs_read_arr(226)(REG_TRIGGER_OH8_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(8 * 9 + 8);
    regs_read_arr(227)(REG_TRIGGER_OH8_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(8 * 9 + 0);
    regs_read_arr(228)(REG_TRIGGER_OH8_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(8 * 9 + 1);
    regs_read_arr(229)(REG_TRIGGER_OH8_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(8 * 9 + 2);
    regs_read_arr(230)(REG_TRIGGER_OH8_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(8 * 9 + 3);
    regs_read_arr(231)(REG_TRIGGER_OH8_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(8 * 9 + 4);
    regs_read_arr(232)(REG_TRIGGER_OH8_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(8 * 9 + 5);
    regs_read_arr(233)(REG_TRIGGER_OH8_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(8 * 9 + 6);
    regs_read_arr(234)(REG_TRIGGER_OH8_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(8 * 9 + 7);
    regs_read_arr(235)(REG_TRIGGER_OH8_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH8_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(8 * 9 + 8);
    regs_read_arr(236)(REG_TRIGGER_OH8_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH8_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(8)(15 downto 0);
    regs_read_arr(236)(REG_TRIGGER_OH8_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH8_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(8)(31 downto 16);
    regs_read_arr(237)(REG_TRIGGER_OH8_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH8_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(8)(15 downto 0);
    regs_read_arr(237)(REG_TRIGGER_OH8_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH8_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(8)(31 downto 16);
    regs_read_arr(238)(REG_TRIGGER_OH8_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH8_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(8)(15 downto 0);
    regs_read_arr(238)(REG_TRIGGER_OH8_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH8_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(8)(31 downto 16);
    regs_read_arr(239)(REG_TRIGGER_OH8_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH8_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(8)(15 downto 0);
    regs_read_arr(239)(REG_TRIGGER_OH8_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH8_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(8)(31 downto 16);
    regs_read_arr(240)(REG_TRIGGER_OH8_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH8_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(8)(15 downto 0);
    regs_read_arr(240)(REG_TRIGGER_OH8_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH8_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(8)(31 downto 16);
    regs_read_arr(241)(REG_TRIGGER_OH9_TRIGGER_RATE_MSB downto REG_TRIGGER_OH9_TRIGGER_RATE_LSB) <= trigger_rate(9);
    regs_read_arr(242)(REG_TRIGGER_OH9_TRIGGER_CNT_MSB downto REG_TRIGGER_OH9_TRIGGER_CNT_LSB) <= trigger_cnt(9);
    regs_read_arr(243)(REG_TRIGGER_OH9_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 0);
    regs_read_arr(244)(REG_TRIGGER_OH9_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 1);
    regs_read_arr(245)(REG_TRIGGER_OH9_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 2);
    regs_read_arr(246)(REG_TRIGGER_OH9_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 3);
    regs_read_arr(247)(REG_TRIGGER_OH9_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 4);
    regs_read_arr(248)(REG_TRIGGER_OH9_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 5);
    regs_read_arr(249)(REG_TRIGGER_OH9_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 6);
    regs_read_arr(250)(REG_TRIGGER_OH9_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 7);
    regs_read_arr(251)(REG_TRIGGER_OH9_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(9 * 9 + 8);
    regs_read_arr(252)(REG_TRIGGER_OH9_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(9 * 9 + 0);
    regs_read_arr(253)(REG_TRIGGER_OH9_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(9 * 9 + 1);
    regs_read_arr(254)(REG_TRIGGER_OH9_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(9 * 9 + 2);
    regs_read_arr(255)(REG_TRIGGER_OH9_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(9 * 9 + 3);
    regs_read_arr(256)(REG_TRIGGER_OH9_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(9 * 9 + 4);
    regs_read_arr(257)(REG_TRIGGER_OH9_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(9 * 9 + 5);
    regs_read_arr(258)(REG_TRIGGER_OH9_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(9 * 9 + 6);
    regs_read_arr(259)(REG_TRIGGER_OH9_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(9 * 9 + 7);
    regs_read_arr(260)(REG_TRIGGER_OH9_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH9_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(9 * 9 + 8);
    regs_read_arr(261)(REG_TRIGGER_OH9_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH9_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(9)(15 downto 0);
    regs_read_arr(261)(REG_TRIGGER_OH9_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH9_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(9)(31 downto 16);
    regs_read_arr(262)(REG_TRIGGER_OH9_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH9_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(9)(15 downto 0);
    regs_read_arr(262)(REG_TRIGGER_OH9_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH9_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(9)(31 downto 16);
    regs_read_arr(263)(REG_TRIGGER_OH9_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH9_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(9)(15 downto 0);
    regs_read_arr(263)(REG_TRIGGER_OH9_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH9_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(9)(31 downto 16);
    regs_read_arr(264)(REG_TRIGGER_OH9_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH9_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(9)(15 downto 0);
    regs_read_arr(264)(REG_TRIGGER_OH9_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH9_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(9)(31 downto 16);
    regs_read_arr(265)(REG_TRIGGER_OH9_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH9_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(9)(15 downto 0);
    regs_read_arr(265)(REG_TRIGGER_OH9_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH9_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(9)(31 downto 16);
    regs_read_arr(266)(REG_TRIGGER_OH10_TRIGGER_RATE_MSB downto REG_TRIGGER_OH10_TRIGGER_RATE_LSB) <= trigger_rate(10);
    regs_read_arr(267)(REG_TRIGGER_OH10_TRIGGER_CNT_MSB downto REG_TRIGGER_OH10_TRIGGER_CNT_LSB) <= trigger_cnt(10);
    regs_read_arr(268)(REG_TRIGGER_OH10_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 0);
    regs_read_arr(269)(REG_TRIGGER_OH10_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 1);
    regs_read_arr(270)(REG_TRIGGER_OH10_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 2);
    regs_read_arr(271)(REG_TRIGGER_OH10_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 3);
    regs_read_arr(272)(REG_TRIGGER_OH10_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 4);
    regs_read_arr(273)(REG_TRIGGER_OH10_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 5);
    regs_read_arr(274)(REG_TRIGGER_OH10_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 6);
    regs_read_arr(275)(REG_TRIGGER_OH10_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 7);
    regs_read_arr(276)(REG_TRIGGER_OH10_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(10 * 9 + 8);
    regs_read_arr(277)(REG_TRIGGER_OH10_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(10 * 9 + 0);
    regs_read_arr(278)(REG_TRIGGER_OH10_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(10 * 9 + 1);
    regs_read_arr(279)(REG_TRIGGER_OH10_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(10 * 9 + 2);
    regs_read_arr(280)(REG_TRIGGER_OH10_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(10 * 9 + 3);
    regs_read_arr(281)(REG_TRIGGER_OH10_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(10 * 9 + 4);
    regs_read_arr(282)(REG_TRIGGER_OH10_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(10 * 9 + 5);
    regs_read_arr(283)(REG_TRIGGER_OH10_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(10 * 9 + 6);
    regs_read_arr(284)(REG_TRIGGER_OH10_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(10 * 9 + 7);
    regs_read_arr(285)(REG_TRIGGER_OH10_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH10_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(10 * 9 + 8);
    regs_read_arr(286)(REG_TRIGGER_OH10_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH10_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(10)(15 downto 0);
    regs_read_arr(286)(REG_TRIGGER_OH10_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH10_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(10)(31 downto 16);
    regs_read_arr(287)(REG_TRIGGER_OH10_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH10_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(10)(15 downto 0);
    regs_read_arr(287)(REG_TRIGGER_OH10_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH10_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(10)(31 downto 16);
    regs_read_arr(288)(REG_TRIGGER_OH10_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH10_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(10)(15 downto 0);
    regs_read_arr(288)(REG_TRIGGER_OH10_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH10_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(10)(31 downto 16);
    regs_read_arr(289)(REG_TRIGGER_OH10_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH10_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(10)(15 downto 0);
    regs_read_arr(289)(REG_TRIGGER_OH10_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH10_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(10)(31 downto 16);
    regs_read_arr(290)(REG_TRIGGER_OH10_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH10_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(10)(15 downto 0);
    regs_read_arr(290)(REG_TRIGGER_OH10_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH10_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(10)(31 downto 16);
    regs_read_arr(291)(REG_TRIGGER_OH11_TRIGGER_RATE_MSB downto REG_TRIGGER_OH11_TRIGGER_RATE_LSB) <= trigger_rate(11);
    regs_read_arr(292)(REG_TRIGGER_OH11_TRIGGER_CNT_MSB downto REG_TRIGGER_OH11_TRIGGER_CNT_LSB) <= trigger_cnt(11);
    regs_read_arr(293)(REG_TRIGGER_OH11_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 0);
    regs_read_arr(294)(REG_TRIGGER_OH11_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 1);
    regs_read_arr(295)(REG_TRIGGER_OH11_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 2);
    regs_read_arr(296)(REG_TRIGGER_OH11_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 3);
    regs_read_arr(297)(REG_TRIGGER_OH11_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 4);
    regs_read_arr(298)(REG_TRIGGER_OH11_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 5);
    regs_read_arr(299)(REG_TRIGGER_OH11_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 6);
    regs_read_arr(300)(REG_TRIGGER_OH11_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 7);
    regs_read_arr(301)(REG_TRIGGER_OH11_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(11 * 9 + 8);
    regs_read_arr(302)(REG_TRIGGER_OH11_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(11 * 9 + 0);
    regs_read_arr(303)(REG_TRIGGER_OH11_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(11 * 9 + 1);
    regs_read_arr(304)(REG_TRIGGER_OH11_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(11 * 9 + 2);
    regs_read_arr(305)(REG_TRIGGER_OH11_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(11 * 9 + 3);
    regs_read_arr(306)(REG_TRIGGER_OH11_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(11 * 9 + 4);
    regs_read_arr(307)(REG_TRIGGER_OH11_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(11 * 9 + 5);
    regs_read_arr(308)(REG_TRIGGER_OH11_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(11 * 9 + 6);
    regs_read_arr(309)(REG_TRIGGER_OH11_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(11 * 9 + 7);
    regs_read_arr(310)(REG_TRIGGER_OH11_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH11_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(11 * 9 + 8);
    regs_read_arr(311)(REG_TRIGGER_OH11_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH11_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(11)(15 downto 0);
    regs_read_arr(311)(REG_TRIGGER_OH11_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH11_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(11)(31 downto 16);
    regs_read_arr(312)(REG_TRIGGER_OH11_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH11_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(11)(15 downto 0);
    regs_read_arr(312)(REG_TRIGGER_OH11_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH11_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(11)(31 downto 16);
    regs_read_arr(313)(REG_TRIGGER_OH11_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH11_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(11)(15 downto 0);
    regs_read_arr(313)(REG_TRIGGER_OH11_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH11_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(11)(31 downto 16);
    regs_read_arr(314)(REG_TRIGGER_OH11_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH11_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(11)(15 downto 0);
    regs_read_arr(314)(REG_TRIGGER_OH11_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH11_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(11)(31 downto 16);
    regs_read_arr(315)(REG_TRIGGER_OH11_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH11_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(11)(15 downto 0);
    regs_read_arr(315)(REG_TRIGGER_OH11_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH11_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(11)(31 downto 16);

    -- Connect write signals
    oh_mask <= regs_write_arr(2)(REG_TRIGGER_CTRL_OH_KILL_MASK_MSB downto REG_TRIGGER_CTRL_OH_KILL_MASK_LSB);
    sector_id <= regs_write_arr(2)(REG_TRIGGER_CTRL_SECTOR_ID_MSB downto REG_TRIGGER_CTRL_SECTOR_ID_LSB);
    sbitmon_link_select <= regs_write_arr(6)(REG_TRIGGER_SBIT_MONITOR_OH_SELECT_MSB downto REG_TRIGGER_SBIT_MONITOR_OH_SELECT_LSB);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);
    reset_cnt <= regs_write_pulse_arr(1);
    sbitmon_reset <= regs_write_pulse_arr(5);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(2)(REG_TRIGGER_CTRL_OH_KILL_MASK_MSB downto REG_TRIGGER_CTRL_OH_KILL_MASK_LSB) <= REG_TRIGGER_CTRL_OH_KILL_MASK_DEFAULT;
    regs_defaults(2)(REG_TRIGGER_CTRL_SECTOR_ID_MSB downto REG_TRIGGER_CTRL_SECTOR_ID_LSB) <= REG_TRIGGER_CTRL_SECTOR_ID_DEFAULT;
    regs_defaults(6)(REG_TRIGGER_SBIT_MONITOR_OH_SELECT_MSB downto REG_TRIGGER_SBIT_MONITOR_OH_SELECT_LSB) <= REG_TRIGGER_SBIT_MONITOR_OH_SELECT_DEFAULT;

    -- Define writable regs
    regs_writable_arr(2) <= '1';
    regs_writable_arr(6) <= '1';

    --==== Registers end ============================================================================
        
end trigger_arch;
