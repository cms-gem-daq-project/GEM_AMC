------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    20:38:00 2016-08-30
-- Module Name:    GEM_TESTS
-- Description:    This module is the entry point for hardware tests e.g. fiber loopback testing with generated data 
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity gem_tests is
    generic(
        g_NUM_OF_OHs        : integer;
        g_NUM_GBTS_PER_OH   : integer;
        g_GEM_STATION       : integer
    );
    port(
        -- reset
        reset_i                     : in  std_logic;
        
        -- TTC
        ttc_clk_i                   : in  t_ttc_clks;        
        ttc_cmds_i                  : in  t_ttc_cmds;
        
        -- Test control
        loopback_gbt_test_en_i      : in std_logic;
        
        -- GBT links
        gbt_link_ready_i            : in  std_logic_vector(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
        gbt_tx_data_arr_o           : out t_gbt_frame_array(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
        gbt_wide_rx_data_arr_i      : in  t_gbt_wide_frame_array(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
        
        -- VFAT3 daq input for channel monitoring
        vfat3_daq_links_arr_i       : in t_oh_vfat_daq_link_arr(g_NUM_OF_OHs - 1 downto 0);
        
        -- IPbus
        ipb_reset_i                 : in  std_logic;
        ipb_clk_i                   : in  std_logic;
        ipb_miso_o                  : out ipb_rbus;
        ipb_mosi_i                  : in  ipb_wbus        
    );
end gem_tests;

architecture Behavioral of gem_tests is

    -- reset
    signal reset_global                 : std_logic;
    signal reset_local                  : std_logic;
    signal reset                        : std_logic;

    -- control
    signal gbt_loop_reset               : std_logic;
    signal gbt_loop_oh_select           : std_logic_vector(3 downto 0);
    signal gbt_loop_err_inject          : std_logic;

    -- gbt loopback oh links
    signal gbt_loop_oh_tx_links_arr     : t_gbt_frame_array(g_NUM_GBTS_PER_OH - 1 downto 0);
    signal gbt_loop_oh_rx_links_arr     : t_gbt_wide_frame_array(g_NUM_GBTS_PER_OH - 1 downto 0);
    
    -- gbt loopback status
    signal gbt_loop_locked_arr          : std_logic_vector(g_NUM_GBTS_PER_OH * 14 - 1 downto 0);
    signal gbt_loop_mega_word_cnt_arr   : t_std32_array(g_NUM_GBTS_PER_OH * 14 - 1 downto 0);
    signal gbt_loop_error_cnt_arr       : t_std32_array(g_NUM_GBTS_PER_OH * 14 - 1 downto 0);
    
    -- VFAT3 DAQ monitor
    signal vfat_daq_links24             : t_vfat_daq_link_arr(23 downto 0);
    signal vfat_daqmon_reset            : std_logic;
    signal vfat_daqmon_enable           : std_logic;
    signal vfat_daqmon_oh_select        : std_logic_vector(3 downto 0);
    signal vfat_daqmon_chan_select      : std_logic_vector(6 downto 0);
    signal vfat_daqmon_chan_global_or   : std_logic;
    signal vfat_daqmon_good_evt_cnt_arr : t_std16_array(23 downto 0); 
    signal vfat_daqmon_chan_fire_cnt_arr: t_std16_array(23 downto 0); 
    
    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------    

begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clk_i.clk_40,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    --== GBT loopback test ==--
    
    g_use_gbtx : if (g_GEM_STATION = 1) or (g_GEM_STATION = 2) generate
        
        -- instantiate the OH tester
        i_oh_prbs_test : entity work.gbt_prbs_loopback_test
            generic map(
                g_NUM_GBTS_PER_OH => g_NUM_GBTS_PER_OH,
                g_TX_ELINKS_PER_GBT  => 10,
                g_RX_ELINKS_PER_GBT  => 14
            )
            port map(
                reset_i                 => reset or gbt_loop_reset,
                enable_i                => loopback_gbt_test_en_i,
                gbt_clk_i               => ttc_clk_i.clk_40,
                gbt_tx_data_arr_o       => gbt_loop_oh_tx_links_arr,
                gbt_wide_rx_data_arr_i  => gbt_loop_oh_rx_links_arr,
                error_inject_en_i       => gbt_loop_err_inject,
                elink_prbs_locked_arr_o => gbt_loop_locked_arr,
                elink_mwords_cnt_arr_o  => gbt_loop_mega_word_cnt_arr,
                elink_error_cnt_arr_o   => gbt_loop_error_cnt_arr
            );
        
        -- fanout the tester TX to all OHs
        g_tx_ohs : for oh in 0 to g_NUM_OF_OHs - 1 generate
            g_tx_gbt : for gbt in 0 to g_NUM_GBTS_PER_OH - 1 generate
                gbt_tx_data_arr_o(oh * g_NUM_GBTS_PER_OH + gbt) <= gbt_loop_oh_tx_links_arr(gbt);
            end generate;
        end generate;
        
        -- MUX the gbt RX links, and route the selected OH to the tester
        g_rx_gbt : for gbt in 0 to g_NUM_GBTS_PER_OH - 1 generate
            gbt_loop_oh_rx_links_arr(gbt) <= gbt_wide_rx_data_arr_i(to_integer(unsigned(gbt_loop_oh_select)) * g_NUM_GBTS_PER_OH + gbt);
        end generate;
        
    end generate;

    --== VFAT3 DAQ monitor ==--
    
    vfat_daq_links24 <= vfat3_daq_links_arr_i(to_integer(unsigned(vfat_daqmon_oh_select)));
    
    g_vfat3_daq_monitors : for i in 0 to 23 generate
        
        i_vfat3_daq_monitor : entity work.vfat3_daq_monitor
            port map(
                reset_i           => reset or vfat_daqmon_reset,
                enable_i          => vfat_daqmon_enable,
                ttc_clk_i         => ttc_clk_i,
                data_en_i         => vfat_daq_links24(i).data_en,
                data_i            => vfat_daq_links24(i).data,
                event_done_i      => vfat_daq_links24(i).event_done,
                crc_error_i       => vfat_daq_links24(i).crc_error,
                chan_global_or_i  => vfat_daqmon_chan_global_or,
                chan_single_idx_i => vfat_daqmon_chan_select,
                cnt_good_events_o => vfat_daqmon_good_evt_cnt_arr(i),
                cnt_chan_fired_o  => vfat_daqmon_chan_fire_cnt_arr(i)
            );
        
    end generate; 
    
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_GEM_TESTS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_GEM_TESTS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_GEM_TESTS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => ttc_clk_i.clk_40,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0000";
    regs_addresses(1)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1000";
    regs_addresses(2)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1001";
    regs_addresses(3)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1002";
    regs_addresses(4)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1010";
    regs_addresses(5)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1011";
    regs_addresses(6)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1012";
    regs_addresses(7)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1013";
    regs_addresses(8)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1014";
    regs_addresses(9)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1015";
    regs_addresses(10)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1016";
    regs_addresses(11)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1017";
    regs_addresses(12)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1018";
    regs_addresses(13)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1019";
    regs_addresses(14)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"101a";
    regs_addresses(15)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"101b";
    regs_addresses(16)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"101c";
    regs_addresses(17)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"101d";
    regs_addresses(18)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"101e";
    regs_addresses(19)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"101f";
    regs_addresses(20)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1020";
    regs_addresses(21)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1021";
    regs_addresses(22)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1022";
    regs_addresses(23)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1023";
    regs_addresses(24)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1024";
    regs_addresses(25)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1025";
    regs_addresses(26)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1026";
    regs_addresses(27)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1027";
    regs_addresses(28)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1028";
    regs_addresses(29)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1029";
    regs_addresses(30)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"102a";
    regs_addresses(31)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"102b";
    regs_addresses(32)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1110";
    regs_addresses(33)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1111";
    regs_addresses(34)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1112";
    regs_addresses(35)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1113";
    regs_addresses(36)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1114";
    regs_addresses(37)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1115";
    regs_addresses(38)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1116";
    regs_addresses(39)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1117";
    regs_addresses(40)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1118";
    regs_addresses(41)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1119";
    regs_addresses(42)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"111a";
    regs_addresses(43)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"111b";
    regs_addresses(44)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"111c";
    regs_addresses(45)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"111d";
    regs_addresses(46)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"111e";
    regs_addresses(47)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"111f";
    regs_addresses(48)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1120";
    regs_addresses(49)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1121";
    regs_addresses(50)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1122";
    regs_addresses(51)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1123";
    regs_addresses(52)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1124";
    regs_addresses(53)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1125";
    regs_addresses(54)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1126";
    regs_addresses(55)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1127";
    regs_addresses(56)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1128";
    regs_addresses(57)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1129";
    regs_addresses(58)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"112a";
    regs_addresses(59)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"112b";
    regs_addresses(60)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1210";
    regs_addresses(61)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1211";
    regs_addresses(62)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1212";
    regs_addresses(63)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1213";
    regs_addresses(64)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1214";
    regs_addresses(65)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1215";
    regs_addresses(66)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1216";
    regs_addresses(67)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1217";
    regs_addresses(68)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1218";
    regs_addresses(69)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1219";
    regs_addresses(70)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"121a";
    regs_addresses(71)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"121b";
    regs_addresses(72)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"121c";
    regs_addresses(73)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"121d";
    regs_addresses(74)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"121e";
    regs_addresses(75)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"121f";
    regs_addresses(76)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1220";
    regs_addresses(77)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1221";
    regs_addresses(78)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1222";
    regs_addresses(79)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1223";
    regs_addresses(80)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1224";
    regs_addresses(81)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1225";
    regs_addresses(82)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1226";
    regs_addresses(83)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1227";
    regs_addresses(84)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1228";
    regs_addresses(85)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1229";
    regs_addresses(86)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"122a";
    regs_addresses(87)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"122b";
    regs_addresses(88)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2000";
    regs_addresses(89)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2001";
    regs_addresses(90)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2010";
    regs_addresses(91)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2020";
    regs_addresses(92)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2030";
    regs_addresses(93)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2040";
    regs_addresses(94)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2050";
    regs_addresses(95)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2060";
    regs_addresses(96)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2070";
    regs_addresses(97)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2080";
    regs_addresses(98)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2090";
    regs_addresses(99)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20a0";
    regs_addresses(100)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20b0";
    regs_addresses(101)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20c0";
    regs_addresses(102)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20d0";
    regs_addresses(103)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20e0";
    regs_addresses(104)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20f0";
    regs_addresses(105)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2100";
    regs_addresses(106)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2110";
    regs_addresses(107)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2120";
    regs_addresses(108)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2130";
    regs_addresses(109)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2140";
    regs_addresses(110)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2150";
    regs_addresses(111)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2160";
    regs_addresses(112)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2170";
    regs_addresses(113)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2180";

    -- Connect read signals
    regs_read_arr(2)(REG_GEM_TESTS_OH_LOOPBACK_CTRL_OH_SELECT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_CTRL_OH_SELECT_LSB) <= gbt_loop_oh_select;
    regs_read_arr(4)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_0_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_0_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 0)(30 downto 0);
    regs_read_arr(4)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_0_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 0);
    regs_read_arr(5)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_0_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 0);
    regs_read_arr(6)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_1_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_1_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 1)(30 downto 0);
    regs_read_arr(6)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_1_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 1);
    regs_read_arr(7)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_1_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 1);
    regs_read_arr(8)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_2_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_2_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 2)(30 downto 0);
    regs_read_arr(8)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_2_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 2);
    regs_read_arr(9)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_2_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_2_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 2);
    regs_read_arr(10)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_3_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_3_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 3)(30 downto 0);
    regs_read_arr(10)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_3_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 3);
    regs_read_arr(11)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_3_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_3_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 3);
    regs_read_arr(12)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_4_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_4_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 4)(30 downto 0);
    regs_read_arr(12)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_4_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 4);
    regs_read_arr(13)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_4_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_4_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 4);
    regs_read_arr(14)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_5_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_5_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 5)(30 downto 0);
    regs_read_arr(14)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_5_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 5);
    regs_read_arr(15)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_5_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_5_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 5);
    regs_read_arr(16)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_6_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_6_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 6)(30 downto 0);
    regs_read_arr(16)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_6_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 6);
    regs_read_arr(17)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_6_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_6_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 6);
    regs_read_arr(18)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_7_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_7_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 7)(30 downto 0);
    regs_read_arr(18)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_7_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 7);
    regs_read_arr(19)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_7_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_7_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 7);
    regs_read_arr(20)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_8_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_8_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 8)(30 downto 0);
    regs_read_arr(20)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_8_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 8);
    regs_read_arr(21)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_8_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_8_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 8);
    regs_read_arr(22)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_9_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_9_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 9)(30 downto 0);
    regs_read_arr(22)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_9_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 9);
    regs_read_arr(23)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_9_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_9_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 9);
    regs_read_arr(24)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_10_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_10_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 10)(30 downto 0);
    regs_read_arr(24)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_10_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 10);
    regs_read_arr(25)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_10_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_10_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 10);
    regs_read_arr(26)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_11_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_11_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 11)(30 downto 0);
    regs_read_arr(26)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_11_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 11);
    regs_read_arr(27)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_11_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_11_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 11);
    regs_read_arr(28)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_12_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_12_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 12)(30 downto 0);
    regs_read_arr(28)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_12_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 12);
    regs_read_arr(29)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_12_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_12_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 12);
    regs_read_arr(30)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_13_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_13_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0 * 14 + 13)(30 downto 0);
    regs_read_arr(30)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_13_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(0 * 14 + 13);
    regs_read_arr(31)(REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_13_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_0_ELINK_13_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0 * 14 + 13);
    regs_read_arr(32)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_0_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_0_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 0)(30 downto 0);
    regs_read_arr(32)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_0_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 0);
    regs_read_arr(33)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_0_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 0);
    regs_read_arr(34)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_1_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_1_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 1)(30 downto 0);
    regs_read_arr(34)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_1_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 1);
    regs_read_arr(35)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_1_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 1);
    regs_read_arr(36)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_2_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_2_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 2)(30 downto 0);
    regs_read_arr(36)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_2_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 2);
    regs_read_arr(37)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_2_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_2_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 2);
    regs_read_arr(38)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_3_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_3_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 3)(30 downto 0);
    regs_read_arr(38)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_3_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 3);
    regs_read_arr(39)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_3_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_3_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 3);
    regs_read_arr(40)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_4_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_4_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 4)(30 downto 0);
    regs_read_arr(40)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_4_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 4);
    regs_read_arr(41)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_4_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_4_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 4);
    regs_read_arr(42)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_5_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_5_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 5)(30 downto 0);
    regs_read_arr(42)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_5_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 5);
    regs_read_arr(43)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_5_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_5_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 5);
    regs_read_arr(44)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_6_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_6_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 6)(30 downto 0);
    regs_read_arr(44)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_6_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 6);
    regs_read_arr(45)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_6_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_6_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 6);
    regs_read_arr(46)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_7_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_7_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 7)(30 downto 0);
    regs_read_arr(46)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_7_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 7);
    regs_read_arr(47)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_7_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_7_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 7);
    regs_read_arr(48)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_8_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_8_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 8)(30 downto 0);
    regs_read_arr(48)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_8_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 8);
    regs_read_arr(49)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_8_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_8_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 8);
    regs_read_arr(50)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_9_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_9_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 9)(30 downto 0);
    regs_read_arr(50)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_9_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 9);
    regs_read_arr(51)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_9_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_9_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 9);
    regs_read_arr(52)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_10_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_10_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 10)(30 downto 0);
    regs_read_arr(52)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_10_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 10);
    regs_read_arr(53)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_10_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_10_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 10);
    regs_read_arr(54)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_11_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_11_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 11)(30 downto 0);
    regs_read_arr(54)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_11_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 11);
    regs_read_arr(55)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_11_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_11_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 11);
    regs_read_arr(56)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_12_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_12_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 12)(30 downto 0);
    regs_read_arr(56)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_12_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 12);
    regs_read_arr(57)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_12_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_12_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 12);
    regs_read_arr(58)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_13_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_13_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1 * 14 + 13)(30 downto 0);
    regs_read_arr(58)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_13_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(1 * 14 + 13);
    regs_read_arr(59)(REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_13_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_1_ELINK_13_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1 * 14 + 13);
    regs_read_arr(60)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_0_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_0_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 0)(30 downto 0);
    regs_read_arr(60)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_0_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 0);
    regs_read_arr(61)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_0_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 0);
    regs_read_arr(62)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_1_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_1_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 1)(30 downto 0);
    regs_read_arr(62)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_1_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 1);
    regs_read_arr(63)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_1_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 1);
    regs_read_arr(64)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_2_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_2_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 2)(30 downto 0);
    regs_read_arr(64)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_2_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 2);
    regs_read_arr(65)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_2_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_2_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 2);
    regs_read_arr(66)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_3_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_3_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 3)(30 downto 0);
    regs_read_arr(66)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_3_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 3);
    regs_read_arr(67)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_3_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_3_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 3);
    regs_read_arr(68)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_4_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_4_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 4)(30 downto 0);
    regs_read_arr(68)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_4_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 4);
    regs_read_arr(69)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_4_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_4_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 4);
    regs_read_arr(70)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_5_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_5_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 5)(30 downto 0);
    regs_read_arr(70)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_5_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 5);
    regs_read_arr(71)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_5_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_5_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 5);
    regs_read_arr(72)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_6_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_6_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 6)(30 downto 0);
    regs_read_arr(72)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_6_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 6);
    regs_read_arr(73)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_6_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_6_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 6);
    regs_read_arr(74)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_7_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_7_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 7)(30 downto 0);
    regs_read_arr(74)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_7_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 7);
    regs_read_arr(75)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_7_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_7_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 7);
    regs_read_arr(76)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_8_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_8_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 8)(30 downto 0);
    regs_read_arr(76)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_8_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 8);
    regs_read_arr(77)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_8_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_8_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 8);
    regs_read_arr(78)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_9_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_9_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 9)(30 downto 0);
    regs_read_arr(78)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_9_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 9);
    regs_read_arr(79)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_9_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_9_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 9);
    regs_read_arr(80)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_10_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_10_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 10)(30 downto 0);
    regs_read_arr(80)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_10_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 10);
    regs_read_arr(81)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_10_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_10_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 10);
    regs_read_arr(82)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_11_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_11_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 11)(30 downto 0);
    regs_read_arr(82)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_11_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 11);
    regs_read_arr(83)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_11_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_11_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 11);
    regs_read_arr(84)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_12_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_12_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 12)(30 downto 0);
    regs_read_arr(84)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_12_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 12);
    regs_read_arr(85)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_12_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_12_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 12);
    regs_read_arr(86)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_13_ERROR_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_13_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2 * 14 + 13)(30 downto 0);
    regs_read_arr(86)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_13_PRBS_LOCKED_BIT) <= gbt_loop_locked_arr(2 * 14 + 13);
    regs_read_arr(87)(REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_13_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_GBT_2_ELINK_13_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2 * 14 + 13);
    regs_read_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_ENABLE_BIT) <= vfat_daqmon_enable;
    regs_read_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_OH_SELECT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_OH_SELECT_LSB) <= vfat_daqmon_oh_select;
    regs_read_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_SELECT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_SELECT_LSB) <= vfat_daqmon_chan_select;
    regs_read_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_GLOBAL_OR_BIT) <= vfat_daqmon_chan_global_or;
    regs_read_arr(90)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT0_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT0_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(0);
    regs_read_arr(90)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT0_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT0_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(0);
    regs_read_arr(91)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT1_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT1_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(1);
    regs_read_arr(91)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT1_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT1_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(1);
    regs_read_arr(92)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT2_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT2_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(2);
    regs_read_arr(92)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT2_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT2_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(2);
    regs_read_arr(93)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT3_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT3_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(3);
    regs_read_arr(93)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT3_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT3_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(3);
    regs_read_arr(94)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT4_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT4_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(4);
    regs_read_arr(94)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT4_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT4_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(4);
    regs_read_arr(95)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT5_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT5_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(5);
    regs_read_arr(95)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT5_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT5_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(5);
    regs_read_arr(96)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT6_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT6_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(6);
    regs_read_arr(96)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT6_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT6_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(6);
    regs_read_arr(97)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT7_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT7_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(7);
    regs_read_arr(97)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT7_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT7_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(7);
    regs_read_arr(98)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT8_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT8_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(8);
    regs_read_arr(98)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT8_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT8_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(8);
    regs_read_arr(99)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT9_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT9_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(9);
    regs_read_arr(99)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT9_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT9_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(9);
    regs_read_arr(100)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT10_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT10_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(10);
    regs_read_arr(100)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT10_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT10_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(10);
    regs_read_arr(101)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT11_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT11_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(11);
    regs_read_arr(101)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT11_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT11_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(11);
    regs_read_arr(102)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT12_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT12_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(12);
    regs_read_arr(102)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT12_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT12_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(12);
    regs_read_arr(103)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT13_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT13_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(13);
    regs_read_arr(103)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT13_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT13_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(13);
    regs_read_arr(104)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT14_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT14_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(14);
    regs_read_arr(104)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT14_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT14_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(14);
    regs_read_arr(105)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT15_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT15_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(15);
    regs_read_arr(105)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT15_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT15_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(15);
    regs_read_arr(106)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT16_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT16_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(16);
    regs_read_arr(106)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT16_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT16_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(16);
    regs_read_arr(107)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT17_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT17_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(17);
    regs_read_arr(107)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT17_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT17_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(17);
    regs_read_arr(108)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT18_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT18_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(18);
    regs_read_arr(108)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT18_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT18_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(18);
    regs_read_arr(109)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT19_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT19_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(19);
    regs_read_arr(109)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT19_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT19_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(19);
    regs_read_arr(110)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT20_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT20_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(20);
    regs_read_arr(110)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT20_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT20_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(20);
    regs_read_arr(111)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT21_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT21_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(21);
    regs_read_arr(111)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT21_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT21_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(21);
    regs_read_arr(112)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT22_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT22_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(22);
    regs_read_arr(112)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT22_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT22_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(22);
    regs_read_arr(113)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT23_GOOD_EVENTS_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT23_GOOD_EVENTS_COUNT_LSB) <= vfat_daqmon_good_evt_cnt_arr(23);
    regs_read_arr(113)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT23_CHANNEL_FIRE_COUNT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_VFAT23_CHANNEL_FIRE_COUNT_LSB) <= vfat_daqmon_chan_fire_cnt_arr(23);

    -- Connect write signals
    gbt_loop_oh_select <= regs_write_arr(2)(REG_GEM_TESTS_OH_LOOPBACK_CTRL_OH_SELECT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_CTRL_OH_SELECT_LSB);
    vfat_daqmon_enable <= regs_write_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_ENABLE_BIT);
    vfat_daqmon_oh_select <= regs_write_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_OH_SELECT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_OH_SELECT_LSB);
    vfat_daqmon_chan_select <= regs_write_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_SELECT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_SELECT_LSB);
    vfat_daqmon_chan_global_or <= regs_write_arr(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_GLOBAL_OR_BIT);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);
    gbt_loop_reset <= regs_write_pulse_arr(1);
    gbt_loop_err_inject <= regs_write_pulse_arr(3);
    vfat_daqmon_reset <= regs_write_pulse_arr(88);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(2)(REG_GEM_TESTS_OH_LOOPBACK_CTRL_OH_SELECT_MSB downto REG_GEM_TESTS_OH_LOOPBACK_CTRL_OH_SELECT_LSB) <= REG_GEM_TESTS_OH_LOOPBACK_CTRL_OH_SELECT_DEFAULT;
    regs_defaults(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_ENABLE_BIT) <= REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_ENABLE_DEFAULT;
    regs_defaults(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_OH_SELECT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_OH_SELECT_LSB) <= REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_OH_SELECT_DEFAULT;
    regs_defaults(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_SELECT_MSB downto REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_SELECT_LSB) <= REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_SELECT_DEFAULT;
    regs_defaults(89)(REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_GLOBAL_OR_BIT) <= REG_GEM_TESTS_VFAT_DAQ_MONITOR_CTRL_VFAT_CHANNEL_GLOBAL_OR_DEFAULT;

    -- Define writable regs
    regs_writable_arr(2) <= '1';
    regs_writable_arr(89) <= '1';

    --==== Registers end ============================================================================

end Behavioral;
